--  SMESH SMESHDS : management of mesh data and SMESH document
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMESHDS_SubMesh.cdl
--  Author : Yves FRICAUD, OCC
--  Module : SMESH

class SubMesh from SMESHDS inherits TShared from MMgt

uses 
	Mesh              from SMDS,
	MeshElement       from SMDS,
	MeshNode          from SMDS,
	ListOfInteger     from TColStd,	
	MapOfMeshElement  from SMDS	

is

	Create (M : Mesh from SMDS) returns mutable SubMesh from SMESHDS;
	
	-- Build

	AddElement   (me : mutable; ME : MeshElement from SMDS);

        RemoveElement    (me: mutable; ME : MeshElement from SMDS);

	AddNode    (me : mutable; ME : MeshNode from SMDS);

        RemoveNode (me: mutable; ME : MeshNode from SMDS);

	
	-- Querry

	NbElements (me: mutable) returns Integer from Standard;

	GetElements (me: mutable ) returns MapOfMeshElement from SMDS;
	---C++ : return const &

	GetIDElements (me: mutable) returns ListOfInteger from TColStd;
	---C++ : return const &

	NbNodes (me: mutable) returns Integer from Standard;

	GetNodes (me: mutable ) returns MapOfMeshElement from SMDS;
	---C++ : return const &

	GetIDNodes (me: mutable) returns ListOfInteger from TColStd;
	---C++ : return const &

fields

	myMesh                  : Mesh              from SMDS;
	myElements              : MapOfMeshElement  from SMDS;
	myNodes                 : MapOfMeshElement  from SMDS;

	myListOfEltIDIsUpdate   : Boolean           from Standard;
	myListOfEltID           : ListOfInteger     from TColStd;

	myListOfNodeIDIsUpdate  : Boolean           from Standard;
	myListOfNodeID          : ListOfInteger     from TColStd;
	

end SubMesh;
