--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org or email : webmaster@opencascade.org 
--
--
--
--  File   : SMDSControl.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

package SMDSControl 

	---Purpose: provides classes for controlling the mesh
	--          according to several criteria

uses

    SMDS
    
is

    ---Category: Classes
    --           

    deferred class MeshBoundary;
	class BoundaryEdges;
    
    	class BoundaryFaces;
    
    ---Category: Package methods
    --           
    
    ComputeNeighborFaces(M:Mesh from SMDS; ME: MeshElement from SMDS; idnode1,idnode2: Integer)
    returns Integer;

    ComputeNeighborVolumes(M:Mesh from SMDS; ME: MeshElement from SMDS; idnode1,idnode2,idnode3: Integer)
    returns Integer;

    ComputeNeighborVolumes(M:Mesh from SMDS; ME: MeshElement from SMDS; idnode1,idnode2,idnode3,idnode4: Integer)
    returns Integer;

end SMDSControl;
