-- File:	SMDS_MeshFace.cdl
-- Created:	Wed Jan 23 16:16:09 2002
-- Author:	Jean-Michel BOULCOURT
--		<jmb@coulox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002


deferred class MeshFace from SMDS inherits MeshElement from SMDS

	---Purpose: 

uses
    MeshElement from SMDS

is

    Initialize(ID: Integer; NbConnections : Integer) returns mutable MeshFace;
    
    ComputeKey(me: mutable) is deferred;
    ---Purpose: compute the  ID of the face  based on the  id's of its
    --          bounding nodes

    GetKey(me) returns Integer is redefined static;    
    ---C++: inline

    NbEdges(me) returns Integer
    is redefined virtual;

    Print(me; OS: in out OStream) is redefined virtual;

fields
    myKey : Integer is protected;
    
end MeshFace;
