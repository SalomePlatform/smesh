--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_MapOfMeshElement.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class MapOfMeshElement from SMDS inherits ExtendedMap from SMDS

	---Purpose:  Redefinition/definition  of methods of Map from TCollection

uses
    MeshElement from SMDS

raises
    NoSuchObject from Standard

is
    Create(NbBuckets : Integer =1) returns MapOfMeshElement from SMDS;
   ---Purpose: Creates   a Map with  <NbBuckets> buckets. Without
   --          arguments the map is automatically dimensioned.
   ---C++: inline

    Find(me; K : MeshElement) returns MeshElement
	---Level: Public
	---Purpose: Returns  the Item stored  with the Key  <K> in the Map. 
        ---Trigger: An exception is raised when <K> is not in the map.
    raises NoSuchObject from Standard  
	---C++: alias operator()
	---C++: return const &
    is static;
    
    ChangeFind(me : in out; K : MeshElement) returns MeshElement
	---Level: Public
	---Purpose: Returns the  Item stored with  the Key  <K> in the
	-- Map. This Item can be   modified with  the  syntax
	-- aMap(K) = newItem; 
        ---Trigger: An exception is raised when <K> is not in the map.
	---C++: alias operator()
	---C++: return &
    raises NoSuchObject from Standard 
    is static;

    FindID(me; ID : Integer) returns MeshElement
	---Level: Public
	---Purpose: Returns  the Item stored  with the ID in the Map. 
        ---Trigger: An exception is raised when ID is not in the map.
    raises NoSuchObject from Standard  
	---C++: alias operator()
	---C++: return const &
    is static;
    

    ContainsID(me; ID : Integer) returns Boolean
	---Level: Public
	---Purpose: Returns True  if the ID is stored  in the
	-- map <me>.
    is static;
    
end MapOfMeshElement;
