--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_MeshElementsIterator.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

deferred class MeshElementsIterator from SMDS 

	---Purpose: The Iterator objet to iterate on all faces of a mesh
	--          

uses
    Mesh from SMDS,
    MeshElement from SMDS,
    MapIteratorOfExtendedOrientedMap from SMDS

raises
    NoMoreObject,
    NoSuchObject

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~SMDS_MeshElementsIterator(){Delete();}"

    Initialize(me : in out; M      : Mesh from SMDS)
	---Purpose: Reset the Iterator on the faces of mesh <M>.
    is deferred;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current meshface.
	--          
	---C++: inline
    is static;
    
    Next(me : in out)
	---Purpose: Moves to the next face.
    raises
    	NoMoreObject from Standard
    is static;
    
    Value(me) returns MeshElement from SMDS
	---Purpose: Returns the meshface.
    raises
    	NoSuchObject from Standard
	---C++: return const &
	---C++: inline
    is static;


fields
    myCurrentMeshElement        : MeshElement  from SMDS is protected;
    myMapIterator : MapIteratorOfExtendedOrientedMap from SMDS is protected;
    
end MeshElementsIterator;
