--  SMESH SMESHDS : management of mesh data and SMESH document
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMESHDS_Script.cdl
--  Author : Yves FRICAUD, OCC
--  Module : SMESH

class Command from SMESHDS inherits TShared from MMgt

uses 

	Integer        from Standard,
	Real           from Standard,
	CommandType    from SMESHDS,
	ListOfReal     from TColStd,
	ListOfInteger  from TColStd

is

	Create (aType : CommandType from SMESHDS) returns Command from SMESHDS;

	AddNode(me: mutable; NewNodeID : Integer; x,y,z : Real); 
		
    	AddEdge(me: mutable; NewEdgeID : Integer; idnode1, idnode2 : Integer); 

    	AddFace(me: mutable; NewFaceID : Integer; idnode1, idnode2, idnode3 : Integer);

    	AddFace(me: mutable; NewFaceID : Integer; idnode1, idnode2, idnode3, idnode4 : Integer);

    	AddVolume(me: mutable; NewVolID : Integer; idnode1, idnode2, idnode3, idnode4 : Integer);

    	AddVolume(me: mutable; NewVolID : Integer; idnode1, idnode2, idnode3, idnode4, idnode5 : Integer);

    	AddVolume(me: mutable; NewVolID : Integer; idnode1, idnode2, idnode3, idnode4, idnode5, idnode6 : Integer);

    	AddVolume(me: mutable; NewVolID : Integer; idnode1, idnode2, idnode3, idnode4, idnode5, idnode6, idnode7, idnode8 : Integer);
    
	MoveNode(me: mutable; NewNodeID : Integer; x,y,z : Real); 

        RemoveNode (me: mutable; NodeID : Integer);

        RemoveElement(me: mutable; ElementID : Integer);
		
	GetType (me: mutable) returns CommandType from SMESHDS;	
	
	GetNumber (me: mutable) returns Integer from Standard;

	GetIndexes 	(me: mutable) 
	---C++ :return const &		
	returns  ListOfInteger  from TColStd;

	GetCoords 	(me: mutable) 
	---C++ :return const &		
	returns  ListOfReal  from TColStd;



fields
	myType     : CommandType from SMESHDS;	
	myNumber   : Integer from Standard;	
	myReals    : ListOfReal from TColStd;
	myIntegers : ListOfInteger  from TColStd;
end Script;
