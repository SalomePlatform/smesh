--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org or email : webmaster@opencascade.org 
--
--
--
--  File   : SMDSControl_MeshBoundary.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

deferred class MeshBoundary from SMDSControl inherits TShared from MMgt

	---Purpose:  common   interface  for  classes   which  extract
	--          boundaries from a mesh

uses

    Mesh from SMDS

is
    Initialize;
    ---Purpose: Initialize an empty MeshBoundary


    Initialize (M : Mesh from SMDS);
    ---Purpose: Initialize a MeshBoundary.


    Compute(me: mutable) is deferred;
    
    ResultMesh(me: mutable) returns Mesh from SMDS;
    

fields
    myMesh : Mesh from SMDS is protected;
    myBoundaryMesh : Mesh from SMDS is protected;

end MeshBoundary;
