--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_Position.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

deferred class Position from SMDS inherits  TShared from MMgt

	---Purpose: abstract  class to define  the different positions
	--          of a node related to the underlying geometry (CAD model)

uses
    Pnt from gp,
    TypeOfPosition from SMDS
    
is

    Initialize(aShapeId: Integer; 
    	       aType: TypeOfPosition from SMDS = SMDS_TOP_UNSPEC) 
    returns mutable Position;

    Coords(me) returns Pnt from gp is deferred;
    ---Purpose: returns the resulting 3d point to be set
    --          in the MeshNode instance
    --          must be redefined by inherited classes
    
    GetTypeOfPosition(me) returns TypeOfPosition from SMDS;
    ---Purpose: returns the type of position
    --          
    ---C++: inline
    
    SetShapeId(me: mutable; aShapeId: Integer);
    ---Purpose: Sets the ShapeId of the position
    --          
    ---C++: inline

    GetShapeId(me) returns Integer;
    ---Purpose: Returns the ShapeId of the position
    --          
    ---C++: inline


fields

    myShapeId : Integer;
    myType    : TypeOfPosition from SMDS;    
end Position;
