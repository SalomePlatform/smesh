-- File:	SMDS_MeshElementsIterator.cdl
-- Created:	Thu Jan 24 12:00:41 2002
-- Author:	Jean-Michel BOULCOURT
--		<jmb@coulox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002


deferred class MeshElementsIterator from SMDS 

	---Purpose: The Iterator objet to iterate on all faces of a mesh
	--          

uses
    Mesh from SMDS,
    MeshElement from SMDS,
    MapIteratorOfExtendedOrientedMap from SMDS

raises
    NoMoreObject,
    NoSuchObject

is

    Delete(me:out) is virtual;
    ---C++: alias "Standard_EXPORT virtual ~SMDS_MeshElementsIterator(){Delete();}"

    Initialize(me : in out; M      : Mesh from SMDS)
	---Purpose: Reset the Iterator on the faces of mesh <M>.
    is deferred;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current meshface.
	--          
	---C++: inline
    is static;
    
    Next(me : in out)
	---Purpose: Moves to the next face.
    raises
    	NoMoreObject from Standard
    is static;
    
    Value(me) returns MeshElement from SMDS
	---Purpose: Returns the meshface.
    raises
    	NoSuchObject from Standard
	---C++: return const &
	---C++: inline
    is static;


fields
    myCurrentMeshElement        : MeshElement  from SMDS is protected;
    myMapIterator : MapIteratorOfExtendedOrientedMap from SMDS is protected;
    
end MeshElementsIterator;
