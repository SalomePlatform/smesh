--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_SpacePosition.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class SpacePosition from SMDS inherits Position from SMDS

	---Purpose: used to characterize a MeshNode with a 3D point
	--          in space not related to any underlying geometry (CAD)

uses
    Pnt from gp

is

    Create returns mutable SpacePosition;
    ---Purpose: empty constructor. the coords are not set

    Create(x, y, z : Real) returns mutable SpacePosition;
    
    Create(aCoords : Pnt from gp) returns mutable SpacePosition;
    
    Coords(me) returns Pnt from gp is redefined virtual;
    ---Purpose: returns the resulting 3d point to be set
    --          in the MeshNode instance
    
    SetCoords(me: mutable; x, y, z : Real);
    ---C++: inline
    
    SetCoords(me: mutable; aCoords : Pnt from gp);
    ---C++: inline
    
fields
    myCoords : Pnt from gp;
    
end SpacePosition;
