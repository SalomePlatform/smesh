-- File:	IntPoly_PntHasher.cdl
-- Created:	Wed Jan 23 16:15:04 2002
-- Author:	Jean-Michel BOULCOURT
--		<jmb@coulox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002


class PntHasher from SMDS

uses  Pnt from gp

is    HashCode(myclass; Point : Pnt from gp;
                        Upper : Integer)
      returns Integer;
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	--          range 0..Upper.
	---C++: inline
	
      IsEqual(myclass; Point1,Point2 : Pnt from gp)
      returns Boolean;
	---Purpose: Returns True  when the two  keys are the same. Two
	--          same  keys  must   have  the  same  hashcode,  the
	--          contrary is not necessary.
	---C++: inline
	
end PntHasher;
