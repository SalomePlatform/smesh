--  SMESH SMESHDS : management of mesh data and SMESH document
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMESHDS_Document.cdl
--  Author : Yves FRICAUD, OCC
--  Module : SMESH

class Document from SMESHDS inherits TShared from MMgt

uses 
	Integer                                        from Standard,
	Mesh                                           from SMESHDS,	
	PtrHypothesis                                  from SMESHDS,	
	DataMapOfIntegerMesh                           from SMESHDS,
	DataMapOfIntegerPtrHypothesis                  from SMESHDS,
	DataMapIteratorOfDataMapOfIntegerMesh          from SMESHDS,
	DataMapIteratorOfDataMapOfIntegerPtrHypothesis from SMESHDS
is

	Create (UserID : Integer from Standard) returns mutable Document;

	NewMesh (me : mutable) returns Integer from Standard;

	RemoveMesh (me : mutable; MeshID : Integer from Standard);

	GetMesh (me : mutable; MeshID : Integer from Standard) returns Mesh from SMESHDS; 


	AddHypothesis (me : mutable; H : PtrHypothesis from SMESHDS);

	RemoveHypothesis (me : mutable; HypID : Integer from Standard);

	GetHypothesis (me : mutable; HypID : Integer from Standard) returns PtrHypothesis from SMESHDS;

	NbMeshes     (me : mutable) returns Integer from Standard;

	NbHypothesis (me : mutable) returns Integer from Standard;

	-- Iterator on Meshes
	InitMeshesIterator(me : mutable);
        
 	NextMesh (me : mutable);
		
	MoreMesh (me : mutable) returns Boolean from Standard;
	
	CurrentMesh (me : mutable ) returns Mesh from SMESHDS; 

	
	--Iterator on Hypothesis
	InitHypothesisIterator (me : mutable );

	NextHypothesis (me : mutable );

	MoreHypothesis (me : mutable ) returns Boolean from Standard;

	CurrentHypothesis (me : mutable) returns PtrHypothesis from SMESHDS;	

fields
	myUserID     : Integer                       from Standard;	
	myMeshes     : DataMapOfIntegerMesh          from SMESHDS;
	myHypothesis : DataMapOfIntegerPtrHypothesis from SMESHDS;

	myMeshesIt     : DataMapIteratorOfDataMapOfIntegerMesh            from SMESHDS;
	myHypothesisIt : DataMapIteratorOfDataMapOfIntegerPtrHypothesis from SMESHDS;

end Document;

