--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_MeshElement.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

deferred class MeshElement from SMDS inherits MeshObject from SMDS

	---Purpose:  MeshElement  is the  base class  for  all mesh --
	--           elements that  constitutes  a mesh.  The children
	--          classes will include   elements like  Node,  Edge,
	--          Face, and Volume.

uses
   ListOfMeshElement from SMDS,
   HArray1OfDir from TColgp,
   Dir from gp,
   Vec from gp,
   ElementType from SMDSAbs

raises
   OutOfRange from Standard
   
is
    
    Initialize(ID: Integer; NbConnections : Integer;
    	       Type: ElementType from SMDSAbs) 
    returns mutable MeshElement;

    HashCode (me; Upper : Integer) returns Integer is redefined static;
	    ---Purpose: Returns a hashed value denoting <me>. This value is in
	    --         the range 1..<Upper>.
    	    ---C++: inline

    IsSame(me; other : MeshElement) returns Boolean;
	---Purpose: Returns True if two mesh elements are same but not
	--          necessary the same orientation
        ---C++: inline


    IsEqual(me; other : MeshElement) returns Boolean;
	---Purpose:  Returns True if  two mesh  elements are  same and
	--          havesame orientation
	---C++: inline


    IsNodeInElement(me; idnode: Integer) returns Boolean;
    ---Purpose: returns true or false if idnode is in the list of the
    --          direct connections
    ---C++: inline
    
    GetEdgeDefinedByNodes(me; rank: Integer; idnode1, idnode2 : out Integer) is virtual;
    ---Purpose: returns the idnodes of the ith edge (rank) of the face
    --          rank must be comprised between 1 and myNbConnections included.
    
    GetFaceDefinedByNodes(me; rank: Integer; idnode : Address;nb: out Integer) is virtual;
    ---Purpose: returns the idnodes of the ith edge (rank) of the face
    --          rank must be comprised between 1 and myNbConnections included.
    
    GetConnections(me) returns Address 
    is virtual protected;

    GetConnection(me; rank: Integer) returns Integer is virtual;

    AddInverseElement(me:mutable; ME: MeshElement from SMDS) is virtual;

    InverseElements(me) returns ListOfMeshElement is virtual;
    ---C++: return const &
    
    ClearInverseElements(me: mutable) is virtual;
    
    NbNodes(me) returns Integer;
    ---C++: inline

    NbEdges(me) returns Integer
    is virtual;

    NbFaces(me) returns Integer
    is virtual;

    GetID(me) returns Integer;
    ---Purpose: returns identifier of node
    ---C++: inline

    GetKey(me) returns Integer is deferred;
    ---Purpose: returns key for hashcode


    SetNormal(me: mutable; rank: Integer; vx,vy,vz : Real) is virtual;
    ---Purpose: set the rank th normal of the element

    SetNormal(me: mutable; rank: Integer; v : Vec from gp) is virtual;
    ---Purpose: set the rank th normal of the element

    GetNormal(me:mutable; rank: Integer) returns Dir from gp is virtual;
    ---Purpose: get the rank th normal of the element

    Print(me; OS: in out OStream) is virtual;
   ---Purpose: 
    ---C++:  alias  "friend Standard_EXPORT Standard_OStream& operator << (Standard_OStream& OS, const Handle(SMDS_MeshElement)& );"

    GetType(me) returns ElementType from SMDSAbs;
    ---Purpose: return the mesh element type
    ---C++: inline

fields

    myID      : Integer is protected;
    myType    : ElementType from SMDSAbs;
    myNbNodes : Integer is protected;
    myNormals : HArray1OfDir from TColgp is protected; 

end MeshElement;
