--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_MeshQuadrangle.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class MeshQuadrangle from SMDS inherits MeshFace from SMDS

	---Purpose: 

uses
    MeshElement from SMDS

is

    Create (ID,idnode1,idnode2,idnode3,idnode4: Integer) returns mutable MeshQuadrangle;
    	---Purpose: constructor for a quandrangle
    
    ComputeKey(me: mutable) is redefined static;
    ---Purpose: compute the  ID of the face  based on the  id's of its
    --          bounding nodes
    ---C++: inline

    GetEdgeDefinedByNodes(me; rank: Integer; idnode1, idnode2 : out Integer) is redefined static;
    ---Purpose: returns the idnodes of the ith edge (rank) of the face
    --          rank must be comprised between 1 and myNbConnections included.
    ---C++: inline
    
    GetConnections(me) returns Address is redefined static;
    ---C++: inline

    GetConnection(me; rank: Integer) returns Integer is redefined static;
    ---C++: inline

    SetConnections(me: mutable; idnode1,idnode2,idnode3,idnode4: Integer) is private; 


fields
    
    myNodes : Integer [4];

end MeshQuadrangle;
