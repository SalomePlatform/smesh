-- File:	SMDS_MeshGroup.cdl
-- Created:	Mon Jun  3 11:49:08 2002
-- Author:	Jean-Michel BOULCOURT
--		<jmb@localhost.localdomain>
---Copyright:	 Matra Datavision 2002


class MeshGroup from SMDS inherits MeshObject from SMDS

	---Purpose: 

uses
    Mesh from SMDS,
    MeshElement from SMDS,
    ElementType from SMDSAbs,
    ListOfMeshGroup from SMDS,
    MapOfMeshElement from SMDS

raises

    NoSuchObject from Standard,
    TypeMismatch from Standard

is

    ---=====================================
    ---Category: public API methods
    --           Group creation and deletion
    --======================================

    Create(aMesh: Mesh from SMDS) returns MeshGroup from SMDS;
    ---Purpose: constructor
	
    AddSubGroup(me: mutable) returns MeshGroup from SMDS;
    ---Purpose:  create a  sub  group.  
    --          uses  a private constructor to create an instance of the
    --          subgroup and attahc it the parent group.
    
    RemoveSubGroup(me: mutable; aGroup: MeshGroup from SMDS)
    returns Boolean
    ---Purpose: remove aGroup from the list of Children
    --          if the subgroup does not belong to this, it returns False
    --          (True otherwise)
    is virtual;
    
    RemoveFromParent(me: mutable)
    returns Boolean
    ---Purpose: remove this from its parent
    --          if this has no parent then it returns False (True otherwise)
    is virtual;
    


    ---=====================================
    ---Category: public API methods
    --           Group contents edition
    --======================================

    Clear(me: mutable);
    ---Purpose: clear the group
    --          once the group is cleared, the type is set to All
    --          but the referenced mesh remains.

    Add(me: mutable; ME: MeshElement from SMDS)
    raises TypeMismatch from Standard;
    ---Purpose: add an element to the group

    Remove(me: mutable; ME: MeshElement from SMDS)
    raises NoSuchObject from Standard;
    ---Purpose: remove an element from the group
    --          raises if the element is not in the group

    ---=====================================
    ---Category: public API methods
    --           Group contents exploration
    --======================================

    IsEmpty(me)
    returns Boolean from Standard;
    ---Purpose: check if the group is empty

    Extent(me) returns Integer from Standard;
    ---Purpose: return numner of elements in the group

    Type(me) returns ElementType from SMDSAbs;
    ---Purpose: return current element type
    --          if the group is empty, returns All

    Contains(me; ME : MeshElement from SMDS)
    returns Boolean from Standard;
    ---Purpose: check if the group contains the mesh element

    Elements(me) returns MapOfMeshElement from SMDS;
    ---Purpose: check if the group contains the mesh element
    ---C++: return const &
    ---C++: inline
    
    ---===========================================
    ---Category: private or protected API methods
    --           
    --============================================

    Create(parent: MeshGroup) returns mutable MeshGroup
    ---Purpose: constructor used internally to create subgroup
    --          
    is private;
    

fields
    myMesh     : Mesh from SMDS;
    myType     : ElementType from SMDSAbs;
    myElements : MapOfMeshElement from SMDS;
    myParent   : MeshGroup from SMDS;
    myChildren : ListOfMeshGroup from SMDS;
    
end MeshGroup;
