--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_MeshNode.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class MeshNode from SMDS inherits MeshElement from SMDS

	---Purpose: 
uses
  Pnt from gp,
  MeshEdge from SMDS,
  MeshFace from SMDS,
  MeshVolume from SMDS,
  ListOfMeshElement from SMDS,
  Position from SMDS

is

    Create (ID: Integer; x, y, z : Real) returns mutable MeshNode;
    
    Print(me; OS: in out OStream) is redefined static;    

    GetKey(me) returns Integer is redefined static;    
    ---C++: inline

    X(me) returns Real;
    ---C++: inline

    Y(me) returns Real;
    ---C++: inline

    Z(me) returns Real;
    ---C++: inline

    Pnt(me) returns Pnt from gp;
    ---C++: inline

    SetPnt(me: mutable;P: Pnt from gp);
    ---C++: inline

    AddInverseElement(me:mutable; ME: MeshElement from SMDS) is redefined static;
	---C++: inline

    RemoveInverseElement(me:mutable; parent: MeshElement from SMDS);

    InverseElements(me) returns ListOfMeshElement is redefined static;
    ---C++: return const &
    ---C++: inline

    ClearInverseElements(me: mutable) is redefined static;
    ---C++: inline

    SetPosition(me: mutable; aPos: Position from SMDS);

    GetPosition(me) returns Position from SMDS;

fields
    myPnt : Pnt from gp;
    myInverseElements : ListOfMeshElement from SMDS;   
    myPosition : Position from SMDS;
    
end MeshNode;
