--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org or email : webmaster@opencascade.org 
--
--
--
--  File   : SMDSEdit_Transform.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class Transform from SMDSEdit 

	---Purpose: tool to modify  a Mesh or MeshElements by applying
	--          a transformation

uses
  Mesh from SMDS,
  ListOfMeshElement from SMDS,
  Trsf from gp
  
is
    Create (aMesh : Mesh from SMDS; aTrsf: Trsf from gp) 
    returns Transform from SMDSEdit;
    ---Purpose: create a transform tool on a whole mesh

    Create (aMesh : Mesh from SMDS; aListOfME : ListOfMeshElement from SMDS;
    	    aTrsf : Trsf from gp)
    returns Transform from SMDSEdit;
    ---Purpose: create  a transform  tool to be  applied on a  list of
    --          meshelements from the mesh aMesh. MeshElements from the
    --          list that do not belong to the mesh will not be treated

    Perform (me: in out);
    ---Purpose: Perform  the current transformation on the  Mesh or on
    --          the list of meshelements if it is not empty
    
    SetTrsf(me: in out; aTrsf: Trsf from gp);
    ---Purpose: replace the field myTrsf by the one given in argument
    --          This can be used to apply another transformation on a mesh
    --          without creating another instance of SMDSEdit_Transform

    GetTrsf(me) returns Trsf from gp;
    ---Purpose: returns the stored Trsf
     
    
fields
    myMesh     : Mesh from SMDS;
    myTrsf     : Trsf from gp;
    myListOfME : ListOfMeshElement from SMDS;
end Transform;
