--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org or email : webmaster@opencascade.org 
--
--
--
--  File   : SMDSControl_BoundaryEdges.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class BoundaryEdges from SMDSControl inherits MeshBoundary from SMDSControl

	---Purpose: compute  the boudary edges  of a mesh that  is the
	--          edges that are shared  by only one face the result
	--          is a new  mesh created in the same  factory as the
	--          original mesh that contains only edges

uses

    Mesh from SMDS,
    MapOfMeshElement from SMDS
is

    Create(M: Mesh from SMDS) returns BoundaryEdges from SMDSControl;
    
    Compute(me: mutable) is redefined virtual;

fields

    myBoundaryEdges : MapOfMeshElement from SMDS;
    
end BoundaryEdges;
