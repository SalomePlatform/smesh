-- File      : SMESHDS_Document.cdl
-- Created   : 
-- Author    : Yves FRICAUD, OCC
-- Project   : SALOME
-- Copyright : OCC

class Document from SMESHDS inherits TShared from MMgt

uses 
	Integer                                        from Standard,
	Mesh                                           from SMESHDS,	
	PtrHypothesis                                  from SMESHDS,	
	DataMapOfIntegerMesh                           from SMESHDS,
	DataMapOfIntegerPtrHypothesis                  from SMESHDS,
	DataMapIteratorOfDataMapOfIntegerMesh          from SMESHDS,
	DataMapIteratorOfDataMapOfIntegerPtrHypothesis from SMESHDS
is

	Create (UserID : Integer from Standard) returns mutable Document;

	NewMesh (me : mutable) returns Integer from Standard;

	RemoveMesh (me : mutable; MeshID : Integer from Standard);

	GetMesh (me : mutable; MeshID : Integer from Standard) returns Mesh from SMESHDS; 


	AddHypothesis (me : mutable; H : PtrHypothesis from SMESHDS);

	RemoveHypothesis (me : mutable; HypID : Integer from Standard);

	GetHypothesis (me : mutable; HypID : Integer from Standard) returns PtrHypothesis from SMESHDS;

	NbMeshes     (me : mutable) returns Integer from Standard;

	NbHypothesis (me : mutable) returns Integer from Standard;

	-- Iterator on Meshes
	InitMeshesIterator(me : mutable);
        
 	NextMesh (me : mutable);
		
	MoreMesh (me : mutable) returns Boolean from Standard;
	
	CurrentMesh (me : mutable ) returns Mesh from SMESHDS; 

	
	--Iterator on Hypothesis
	InitHypothesisIterator (me : mutable );

	NextHypothesis (me : mutable );

	MoreHypothesis (me : mutable ) returns Boolean from Standard;

	CurrentHypothesis (me : mutable) returns PtrHypothesis from SMESHDS;	

fields
	myUserID     : Integer                       from Standard;	
	myMeshes     : DataMapOfIntegerMesh          from SMESHDS;
	myHypothesis : DataMapOfIntegerPtrHypothesis from SMESHDS;

	myMeshesIt     : DataMapIteratorOfDataMapOfIntegerMesh            from SMESHDS;
	myHypothesisIt : DataMapIteratorOfDataMapOfIntegerPtrHypothesis from SMESHDS;

end Document;

