--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_EdgePosition.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

class EdgePosition from SMDS inherits Position from SMDS

	---Purpose: used to characterize a MeshNode with a CAD edge

uses
    Pnt from gp

is

    Create returns mutable EdgePosition;
    ---Purpose: empty constructor. the edge is not set

    Create(aEdgeId : Integer; aUParam : Real) returns mutable EdgePosition;

    Coords(me) returns Pnt from gp is redefined virtual;
    ---Purpose: returns the resulting 3d point to be set
    --          in the MeshNode instance
    
    SetUParameter(me: mutable; aUparam : Real);
    ---C++: inline

    GetUParameter(me) returns Real;
    ---C++: inline
    
fields

    myUParameter : Real;
    
end EdgePosition;
