--  SMESH SMDS : implementaion of Salome mesh data structure
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMDS_MeshFace.cdl
--  Author : Jean-Michel BOULCOURT
--  Module : SMESH

deferred class MeshFace from SMDS inherits MeshElement from SMDS

	---Purpose: 

uses
    MeshElement from SMDS

is

    Initialize(ID: Integer; NbConnections : Integer) returns mutable MeshFace;
    
    ComputeKey(me: mutable) is deferred;
    ---Purpose: compute the  ID of the face  based on the  id's of its
    --          bounding nodes

    GetKey(me) returns Integer is redefined static;    
    ---C++: inline

    NbEdges(me) returns Integer
    is redefined virtual;

    Print(me; OS: in out OStream) is redefined virtual;

fields
    myKey : Integer is protected;
    
end MeshFace;
