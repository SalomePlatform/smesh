--  SMESH SMESHDS : management of mesh data and SMESH document
--
--  Copyright (C) 2003  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
--  CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS 
-- 
--  This library is free software; you can redistribute it and/or 
--  modify it under the terms of the GNU Lesser General Public 
--  License as published by the Free Software Foundation; either 
--  version 2.1 of the License. 
-- 
--  This library is distributed in the hope that it will be useful, 
--  but WITHOUT ANY WARRANTY; without even the implied warranty of 
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
--  Lesser General Public License for more details. 
-- 
--  You should have received a copy of the GNU Lesser General Public 
--  License along with this library; if not, write to the Free Software 
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA 
-- 
--  See http://www.opencascade.org/SALOME/ or email : webmaster.salome@opencascade.org 
--
--
--
--  File   : SMESHDS.cdl
--  Author : Yves FRICAUD, OCC
--  Module : SMESH

package SMESHDS

uses 
	Standard,
	TColStd,
	SMDS,
	TCollection,
	TopoDS,
	TopTools

is

	enumeration  
	CommandType  is AddNode,  AddEdge,  AddTriangle,  AddQuadrangle,   AddTetrahedron,  AddPyramid,  
	AddPrism,  AddHexahedron, RemoveNode, RemoveElement, MoveNode 
	end CommandType;	
	
	class Document;
	
	class Mesh;

	class SubMesh;

	imported Hypothesis;

	pointer PtrHypothesis to Hypothesis from SMESHDS;
	
	class Script;

	class Command;



	class DataMapOfShapeSubMesh instantiates DataMap from TCollection (Shape from TopoDS,
									   SubMesh from SMESHDS,
								           ShapeMapHasher from TopTools);

	class DataMapOfIntegerSubMesh instantiates  DataMap from TCollection (Integer          from Standard,
								              SubMesh          from SMESHDS,
								              MapIntegerHasher from TColStd);	


	class DataMapOfIntegerPtrHypothesis instantiates  DataMap from TCollection (Integer from Standard,
									            PtrHypothesis from SMESHDS,
										    MapIntegerHasher from TColStd);	
											
	class DataMapOfIntegerMesh instantiates  DataMap from TCollection (Integer from Standard,
								           Mesh    from SMESHDS,
								           MapIntegerHasher from TColStd);	
											    
	class ListOfPtrHypothesis instantiates List from TCollection (PtrHypothesis from SMESHDS);

	
	class DataMapOfShapeListOfPtrHypothesis instantiates DataMap from TCollection (Shape from TopoDS,
								       	    	    ListOfPtrHypothesis from SMESHDS, 
										    ShapeMapHasher from TopTools);

	class ListOfAsciiString  instantiates List from TCollection (AsciiString from TCollection);

	class ListOfCommand      instantiates List from TCollection (Command from SMESHDS);
								 

end SMESHDS;