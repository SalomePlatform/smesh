-- File:	SMDS_MeshNode.cdl
-- Created:	Wed Jan 23 16:15:04 2002
-- Author:	Jean-Michel BOULCOURT
--		<jmb@coulox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 2002


class MeshNode from SMDS inherits MeshElement from SMDS

	---Purpose: 
uses
  Pnt from gp,
  MeshEdge from SMDS,
  MeshFace from SMDS,
  MeshVolume from SMDS,
  ListOfMeshElement from SMDS,
  Position from SMDS

is

    Create (ID: Integer; x, y, z : Real) returns mutable MeshNode;
    
    Print(me; OS: in out OStream) is redefined static;    

    GetKey(me) returns Integer is redefined static;    
    ---C++: inline

    X(me) returns Real;
    ---C++: inline

    Y(me) returns Real;
    ---C++: inline

    Z(me) returns Real;
    ---C++: inline

    Pnt(me) returns Pnt from gp;
    ---C++: inline

    SetPnt(me: mutable;P: Pnt from gp);
    ---C++: inline

    AddInverseElement(me:mutable; ME: MeshElement from SMDS) is redefined static;
	---C++: inline

    RemoveInverseElement(me:mutable; parent: MeshElement from SMDS);

    InverseElements(me) returns ListOfMeshElement is redefined static;
    ---C++: return const &
    ---C++: inline

    ClearInverseElements(me: mutable) is redefined static;
    ---C++: inline

    SetPosition(me: mutable; aPos: Position from SMDS);

    GetPosition(me) returns Position from SMDS;

fields
    myPnt : Pnt from gp;
    myInverseElements : ListOfMeshElement from SMDS;   
    myPosition : Position from SMDS;
    
end MeshNode;
